ENTITY MULTIPLEXADOR4BITS IS 
	PORT(
		Em14B,Em24B,Em34B,Em44B:IN BIT_VECTOR(3 DOWNTO 0);
		Em11B,Em21B,Em31B,Em41B,Em51B,Em61B:IN BIT;
		S01,S11,S21,S31,BLD:IN BIT;
		VetorSaida:OUT BIT_VECTOR(3 DOWNTO 0);
		Cout,Ctrl:OUT BIT);
END MULTIPLEXADOR4BITS;
ARCHITECTURE mux4BIT OF MULTIPLEXADOR4BITS IS
SIGNAL inter:BIT_VECTOR(4 DOWNTO 0);
COMPONENT MULTIPLEXADOR1BIT
PORT(
		Em1,Em2,Em3,Em4,Em5,Em6:IN BIT;
		S0,S1,S2,S3:IN BIT;
		Saida:OUT BIT);
END COMPONENT;
BEGIN
g:FOR i IN 0 TO 3 GENERATE
mux: MULTIPLEXADOR1BIT PORT MAP(Em1=>Em14B(i),Em2=>Em24B(i),Em3=>Em34B(i),Em4=>Em44B(i),Em5=>'0',Em6=>'0',S0=>S01,S1=>S11,S2=>S21,S3=>S31,Saida=>inter(i));
END GENERATE;
muxCout: MULTIPLEXADOR1BIT PORT MAP(Em1=>Em11B,Em2=>Em21B,Em3=>Em31B,Em4=>Em41B,Em5=>Em51B,Em6=>Em61B,S0=>S01,S1=>S11,S2=>S21,S3=>S31,Saida=>inter(4));

VetorSaida(0)<=(BLD) AND inter(0);
VetorSaida(1)<=(BLD) AND inter(1);
VetorSaida(2)<=(BLD) AND inter(2);
VetorSaida(3)<=(BLD) AND inter(3);
Cout<=(BLD) AND inter(4);
Ctrl<= BLD;
END mux4BIT;